add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM1/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM2/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM3/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM4/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM5/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM6/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM7/inst/wea[0]}} 


add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[28]}}


add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[29]}}

add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[30]}}

add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[31]}}


create_debug_core u_ila_0 ila
set_property ALL_PROBE_SAME_MU true [get_debug_cores u_ila_0]
set_property ALL_PROBE_SAME_MU_CNT 4 [get_debug_cores u_ila_0]
set_property C_ADV_TRIGGER true [get_debug_cores u_ila_0]
set_property C_DATA_DEPTH 1024 [get_debug_cores u_ila_0]
set_property C_EN_STRG_QUAL false [get_debug_cores u_ila_0]
set_property C_INPUT_PIPE_STAGES 0 [get_debug_cores u_ila_0]
set_property C_TRIGIN_EN false [get_debug_cores u_ila_0]
set_property C_TRIGOUT_EN false [get_debug_cores u_ila_0]
set_property port_width 1 [get_debug_ports u_ila_0/clk]
connect_debug_port u_ila_0/clk [get_nets [list clk_x3]]
set_property PROBE_TYPE DATA_AND_TRIGGER [get_debug_ports u_ila_0/probe0]
set_property port_width 3 [get_debug_ports u_ila_0/probe0]
connect_debug_port u_ila_0/probe0 [get_nets [list {cpu1/fdem/Pipeline/Load_Store_Op__ex_mem[0]} {cpu1/fdem/Pipeline/Load_Store_Op__ex_mem[1]} {cpu1/fdem/Pipeline/Load_Store_Op__ex_mem[3]}]]
create_debug_port u_ila_0 probe
set_property PROBE_TYPE DATA_AND_TRIGGER [get_debug_ports u_ila_0/probe1]
set_property port_width 32 [get_debug_ports u_ila_0/probe1]
connect_debug_port u_ila_0/probe1 [get_nets [list {cpu1/fdem/Pipeline/PC__IF_ID[0]} {cpu1/fdem/Pipeline/PC__IF_ID[1]} {cpu1/fdem/Pipeline/PC__IF_ID[2]} {cpu1/fdem/Pipeline/PC__IF_ID[3]} {cpu1/fdem/Pipeline/PC__IF_ID[4]} {cpu1/fdem/Pipeline/PC__IF_ID[5]} {cpu1/fdem/Pipeline/PC__IF_ID[6]} {cpu1/fdem/Pipeline/PC__IF_ID[7]} {cpu1/fdem/Pipeline/PC__IF_ID[8]} {cpu1/fdem/Pipeline/PC__IF_ID[9]} {cpu1/fdem/Pipeline/PC__IF_ID[10]} {cpu1/fdem/Pipeline/PC__IF_ID[11]} {cpu1/fdem/Pipeline/PC__IF_ID[12]} {cpu1/fdem/Pipeline/PC__IF_ID[13]} {cpu1/fdem/Pipeline/PC__IF_ID[14]} {cpu1/fdem/Pipeline/PC__IF_ID[15]} {cpu1/fdem/Pipeline/PC__IF_ID[16]} {cpu1/fdem/Pipeline/PC__IF_ID[17]} {cpu1/fdem/Pipeline/PC__IF_ID[18]} {cpu1/fdem/Pipeline/PC__IF_ID[19]} {cpu1/fdem/Pipeline/PC__IF_ID[20]} {cpu1/fdem/Pipeline/PC__IF_ID[21]} {cpu1/fdem/Pipeline/PC__IF_ID[22]} {cpu1/fdem/Pipeline/PC__IF_ID[23]} {cpu1/fdem/Pipeline/PC__IF_ID[24]} {cpu1/fdem/Pipeline/PC__IF_ID[25]} {cpu1/fdem/Pipeline/PC__IF_ID[26]} {cpu1/fdem/Pipeline/PC__IF_ID[27]} {cpu1/fdem/Pipeline/PC__IF_ID[28]} {cpu1/fdem/Pipeline/PC__IF_ID[29]} {cpu1/fdem/Pipeline/PC__IF_ID[30]} {cpu1/fdem/Pipeline/PC__IF_ID[31]}]]
create_debug_port u_ila_0 probe
set_property PROBE_TYPE DATA_AND_TRIGGER [get_debug_ports u_ila_0/probe2]
set_property port_width 32 [get_debug_ports u_ila_0/probe2]
connect_debug_port u_ila_0/probe2 [get_nets [list {cpu1/fdem/Pipeline/proc_addr_port1[0]} {cpu1/fdem/Pipeline/proc_addr_port1[1]} {cpu1/fdem/Pipeline/proc_addr_port1[2]} {cpu1/fdem/Pipeline/proc_addr_port1[3]} {cpu1/fdem/Pipeline/proc_addr_port1[4]} {cpu1/fdem/Pipeline/proc_addr_port1[5]} {cpu1/fdem/Pipeline/proc_addr_port1[6]} {cpu1/fdem/Pipeline/proc_addr_port1[7]} {cpu1/fdem/Pipeline/proc_addr_port1[8]} {cpu1/fdem/Pipeline/proc_addr_port1[9]} {cpu1/fdem/Pipeline/proc_addr_port1[10]} {cpu1/fdem/Pipeline/proc_addr_port1[11]} {cpu1/fdem/Pipeline/proc_addr_port1[12]} {cpu1/fdem/Pipeline/proc_addr_port1[13]} {cpu1/fdem/Pipeline/proc_addr_port1[14]} {cpu1/fdem/Pipeline/proc_addr_port1[15]} {cpu1/fdem/Pipeline/proc_addr_port1[16]} {cpu1/fdem/Pipeline/proc_addr_port1[17]} {cpu1/fdem/Pipeline/proc_addr_port1[18]} {cpu1/fdem/Pipeline/proc_addr_port1[19]} {cpu1/fdem/Pipeline/proc_addr_port1[20]} {cpu1/fdem/Pipeline/proc_addr_port1[21]} {cpu1/fdem/Pipeline/proc_addr_port1[22]} {cpu1/fdem/Pipeline/proc_addr_port1[23]} {cpu1/fdem/Pipeline/proc_addr_port1[24]} {cpu1/fdem/Pipeline/proc_addr_port1[25]} {cpu1/fdem/Pipeline/proc_addr_port1[26]} {cpu1/fdem/Pipeline/proc_addr_port1[27]} {cpu1/fdem/Pipeline/proc_addr_port1[28]} {cpu1/fdem/Pipeline/proc_addr_port1[29]} {cpu1/fdem/Pipeline/proc_addr_port1[30]} {cpu1/fdem/Pipeline/proc_addr_port1[31]}]]
create_debug_port u_ila_0 probe
set_property PROBE_TYPE DATA_AND_TRIGGER [get_debug_ports u_ila_0/probe3]
set_property port_width 32 [get_debug_ports u_ila_0/probe3]
connect_debug_port u_ila_0/probe3 [get_nets [list {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[0]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[1]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[2]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[3]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[4]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[5]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[6]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[7]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[8]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[9]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[10]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[11]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[12]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[13]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[14]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[15]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[16]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[17]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[18]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[19]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[20]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[21]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[22]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[23]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[24]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[25]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[26]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[27]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[28]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[29]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[30]} {cpu1/fdem/Pipeline/VECTOR_UNIT/proc_din[31]}]]
set_property C_CLK_INPUT_FREQ_HZ 300000000 [get_debug_cores dbg_hub]
set_property C_ENABLE_CLK_DIVIDER false [get_debug_cores dbg_hub]
set_property C_USER_SCAN_CHAIN 1 [get_debug_cores dbg_hub]
connect_debug_port dbg_hub/clk [get_nets clk_int]